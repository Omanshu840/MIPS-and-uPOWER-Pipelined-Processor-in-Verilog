module PCmux(Y, D0, D1, S);

    output [63:0] Y;
    input [63:0] D0, D1;
    input S;

    mux21 m1(Y[0], D0[0], D1[0], S);
    mux21 m2(Y[1], D0[1], D1[1], S);
    mux21 m3(Y[2], D0[2], D1[2], S);
    mux21 m4(Y[3], D0[3], D1[3], S);
    mux21 m5(Y[4], D0[4], D1[4], S);
    mux21 m6(Y[5], D0[5], D1[5], S);
    mux21 m7(Y[6], D0[6], D1[6], S);
    mux21 m8(Y[7], D0[7], D1[7], S);
    mux21 m9(Y[8], D0[8], D1[8], S);
    mux21 m10(Y[9], D0[9], D1[9], S);
    mux21 m11(Y[10], D0[10], D1[10], S);
    mux21 m12(Y[11], D0[11], D1[11], S);
    mux21 m13(Y[12], D0[12], D1[12], S);
    mux21 m14(Y[13], D0[13], D1[13], S);
    mux21 m15(Y[14], D0[14], D1[14], S);
    mux21 m16(Y[15], D0[15], D1[15], S);
    mux21 m17(Y[16], D0[16], D1[16], S);
    mux21 m18(Y[17], D0[17], D1[17], S);
    mux21 m19(Y[18], D0[18], D1[18], S);
    mux21 m20(Y[19], D0[19], D1[19], S);
    mux21 m21(Y[20], D0[20], D1[20], S);
    mux21 m22(Y[21], D0[21], D1[21], S);
    mux21 m23(Y[22], D0[22], D1[22], S);
    mux21 m24(Y[23], D0[23], D1[23], S);
    mux21 m25(Y[24], D0[24], D1[24], S);
    mux21 m26(Y[25], D0[25], D1[25], S);
    mux21 m27(Y[26], D0[26], D1[26], S);
    mux21 m28(Y[27], D0[27], D1[27], S);
    mux21 m29(Y[28], D0[28], D1[28], S);
    mux21 m30(Y[29], D0[29], D1[29], S);
    mux21 m31(Y[30], D0[30], D1[30], S);
    mux21 m32(Y[31], D0[31], D1[31], S);
    mux21 m33(Y[32], D0[32], D1[32], S);
    mux21 m34(Y[33], D0[33], D1[33], S);
    mux21 m35(Y[34], D0[34], D1[34], S);
    mux21 m36(Y[35], D0[35], D1[35], S);
    mux21 m37(Y[36], D0[36], D1[36], S);
    mux21 m38(Y[37], D0[37], D1[37], S);
    mux21 m39(Y[38], D0[38], D1[38], S);
    mux21 m40(Y[39], D0[39], D1[39], S);
    mux21 m41(Y[40], D0[40], D1[40], S);
    mux21 m42(Y[41], D0[41], D1[41], S);
    mux21 m43(Y[42], D0[42], D1[42], S);
    mux21 m44(Y[43], D0[43], D1[43], S);
    mux21 m45(Y[44], D0[44], D1[44], S);
    mux21 m46(Y[45], D0[45], D1[45], S);
    mux21 m47(Y[46], D0[46], D1[46], S);
    mux21 m48(Y[47], D0[47], D1[47], S);
    mux21 m49(Y[48], D0[48], D1[48], S);
    mux21 m50(Y[49], D0[49], D1[49], S);
    mux21 m51(Y[50], D0[50], D1[50], S);
    mux21 m52(Y[51], D0[51], D1[51], S);
    mux21 m53(Y[52], D0[52], D1[52], S);
    mux21 m54(Y[53], D0[53], D1[53], S);
    mux21 m55(Y[54], D0[54], D1[54], S);
    mux21 m56(Y[55], D0[55], D1[55], S);
    mux21 m57(Y[56], D0[56], D1[56], S);
    mux21 m58(Y[57], D0[57], D1[57], S);
    mux21 m59(Y[58], D0[58], D1[58], S);
    mux21 m60(Y[59], D0[59], D1[59], S);
    mux21 m61(Y[60], D0[60], D1[60], S);
    mux21 m62(Y[61], D0[61], D1[61], S);
    mux21 m63(Y[62], D0[62], D1[62], S);
    mux21 m64(Y[63], D0[63], D1[63], S);

endmodule